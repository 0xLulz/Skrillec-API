module stresser

